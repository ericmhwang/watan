1
1 5 0 5 0 g c  37  25  30 
0 2 0 0 0 g c  32  44 
10 1 0 0 0 g c  16  40 
0 0 3 0 0 g c  20  27 
0 3 1 10 2 5 3 4 4 7 5 10 6 11 7 3 8 8 9 2 10 6 11 8 12 12 13 5 14 11 15 4 16 6 17 9 18 9 
8
